//====================================================================
// simpleEthernet
// eth_rx.v
// Ethernet RMII receive module
// 12/10/24
//====================================================================

module eth_rx (
  input wire Clk,
  input wire Rst,
  input wire [1:0] Rxd,
  input wire Crs_DV
);

endmodule
