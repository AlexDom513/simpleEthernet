// vim: ts=4 sw=4 expandtab

// THIS IS GENERATED VERILOG CODE.
// https://bues.ch/h/crcgen
// 
// This code is Public Domain.
// Permission to use, copy, modify, and/or distribute this software for any
// purpose with or without fee is hereby granted.
// 
// THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
// WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
// MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR ANY
// SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES WHATSOEVER
// RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN ACTION OF CONTRACT,
// NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF OR IN CONNECTION WITH THE
// USE OR PERFORMANCE OF THIS SOFTWARE.

`ifndef CRC_V_
`define CRC_V_

// CRC polynomial coefficients: x^32 + x^26 + x^23 + x^22 + x^16 + x^12 + x^11 + x^10 + x^8 + x^7 + x^5 + x^4 + x^2 + x + 1
//                              0xEDB88320 (hex)
// CRC width:                   32 bits
// CRC shift direction:         right (little endian)
// Input word width:            2 bits

module crc_gen (
  input           Clk,
  input           Rst,
  input           Crc_En,
  input   [1:0]   Data,
  output  [31:0]  Crc_Out
);

  reg [31:0] lfsr_q;
  wire [31:0] lfsr_c;

  // xor on the output
  assign Crc_Out = lfsr_c ^ 32'hFFFFFFFF;

  assign lfsr_c[0] = lfsr_q[2];
  assign lfsr_c[1] = lfsr_q[3];
  assign lfsr_c[2] = lfsr_q[4];
  assign lfsr_c[3] = lfsr_q[5];
  assign lfsr_c[4] = lfsr_q[0] ^ lfsr_q[6] ^ Data[0];
  assign lfsr_c[5] = lfsr_q[1] ^ lfsr_q[7] ^ Data[1];
  assign lfsr_c[6] = lfsr_q[8];
  assign lfsr_c[7] = lfsr_q[0] ^ lfsr_q[9] ^ Data[0];
  assign lfsr_c[8] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[10] ^ Data[0] ^ Data[1];
  assign lfsr_c[9] = lfsr_q[1] ^ lfsr_q[11] ^ Data[1];
  assign lfsr_c[10] = lfsr_q[12];
  assign lfsr_c[11] = lfsr_q[13];
  assign lfsr_c[12] = lfsr_q[14];
  assign lfsr_c[13] = lfsr_q[15];
  assign lfsr_c[14] = lfsr_q[0] ^ lfsr_q[16] ^ Data[0];
  assign lfsr_c[15] = lfsr_q[1] ^ lfsr_q[17] ^ Data[1];
  assign lfsr_c[16] = lfsr_q[18];
  assign lfsr_c[17] = lfsr_q[19];
  assign lfsr_c[18] = lfsr_q[0] ^ lfsr_q[20] ^ Data[0];
  assign lfsr_c[19] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[21] ^ Data[0] ^ Data[1];
  assign lfsr_c[20] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[22] ^ Data[0] ^ Data[1];
  assign lfsr_c[21] = lfsr_q[1] ^ lfsr_q[23] ^ Data[1];
  assign lfsr_c[22] = lfsr_q[0] ^ lfsr_q[24] ^ Data[0];
  assign lfsr_c[23] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[25] ^ Data[0] ^ Data[1];
  assign lfsr_c[24] = lfsr_q[1] ^ lfsr_q[26] ^ Data[1];
  assign lfsr_c[25] = lfsr_q[0] ^ lfsr_q[27] ^ Data[0];
  assign lfsr_c[26] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[28] ^ Data[0] ^ Data[1];
  assign lfsr_c[27] = lfsr_q[1] ^ lfsr_q[29] ^ Data[1];
  assign lfsr_c[28] = lfsr_q[0] ^ lfsr_q[30] ^ Data[0];
  assign lfsr_c[29] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[31] ^ Data[0] ^ Data[1];
  assign lfsr_c[30] = lfsr_q[0] ^ lfsr_q[1] ^ Data[0] ^ Data[1];
  assign lfsr_c[31] = lfsr_q[1] ^ Data[1];

  always @(posedge Clk)
  begin
    if (Rst)
      lfsr_q <= 32'hFFFFFFFF;
    else begin
      if (Crc_En)
        lfsr_q <= lfsr_c;
      else
        lfsr_q <= lfsr_q;
    end
  end

endmodule

`endif // CRC_V_
