//====================================================================
// simpleEthernet
// eth_tx_ctrl.v
// Ethernet RMII transmit module control
// 12/23/24
//====================================================================

module eth_tx_ctrl (
  input wire      Clk,
  input wire      Rst
);

  //==========================================
  // Constants
  //==========================================

  //==========================================
  // Wires/Registers
  //==========================================

  //==========================================
  // eth_ctrl_fsm
  //==========================================

endmodule
